`timescale 1ns / 1ps

module decoder_3x8(a,d);
input [2:0]a;
output [7:0]d;

assign d[0]=(~a[2])&(~a[1])&(~a[0]);
assign d[1]=(~a[2])&(~a[1])&a[0];
assign d[2]=(~a[2])&a[1]&(~a[0]);
assign d[3]=(~a[2])&a[1]&a[0];
assign d[4]=a[2]&(~a[1])&(~a[0]); 
assign d[5]=a[2]&(~a[1])&a[0];
assign d[6]=a[2]&a[1]&(~a[0]); 
assign d[7]=a[2]&a[1]&a[0];
       
endmodule
