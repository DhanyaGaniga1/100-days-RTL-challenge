`timescale 1ns / 1ps

module half_adder(input a,b,output sum,cout);

and g1(cout,a,b);
xor g2(sum,a,b);

endmodule
